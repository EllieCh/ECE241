module andGate(input a, b, output d);
	assign d = a&&b;
endmodule