// Audio_in.v

// Generated using ACDS version 16.0 211

`timescale 1 ps / 1 ps
module Audio_in (
		input  wire        reg_clk,     //       control_clock.clk
		input  wire        reg_reset,   // control_clock_reset.reset
		input  wire        aes_clk,     //   conduit_aes_audio.export
		input  wire        aes_de,      //                    .export
		input  wire        aes_ws,      //                    .export
		input  wire        aes_data,    //                    .export
		input  wire        aud_clk,     //          dout_clock.clk
		input  wire        reset,       //    dout_clock_reset.reset
		input  wire        aud_ready,   //                dout.ready
		output wire        aud_valid,   //                    .valid
		output wire        aud_sop,     //                    .startofpacket
		output wire        aud_eop,     //                    .endofpacket
		output wire [7:0]  aud_channel, //                    .channel
		output wire [23:0] aud_data,    //                    .data
		input  wire [7:0]  channel0,    //     conduit_control.export
		input  wire [7:0]  channel1,    //                    .export
		output wire [7:0]  fifo_status, //                    .export
		input  wire        fifo_reset   //                    .export
	);

	clocked_audio_input #(
		.G_CAI_FIFO_DEPTH       (4),
		.G_CAI_INCLUDE_CTRL_REG (0)
	) audio_in_inst (
		.reg_clk       (reg_clk),     //       control_clock.clk
		.reg_reset     (reg_reset),   // control_clock_reset.reset
		.aes_clk       (aes_clk),     //   conduit_aes_audio.export
		.aes_de        (aes_de),      //                    .export
		.aes_ws        (aes_ws),      //                    .export
		.aes_data      (aes_data),    //                    .export
		.aud_clk       (aud_clk),     //          dout_clock.clk
		.reset         (reset),       //    dout_clock_reset.reset
		.aud_ready     (aud_ready),   //                dout.ready
		.aud_valid     (aud_valid),   //                    .valid
		.aud_sop       (aud_sop),     //                    .startofpacket
		.aud_eop       (aud_eop),     //                    .endofpacket
		.aud_channel   (aud_channel), //                    .channel
		.aud_data      (aud_data),    //                    .data
		.channel0      (channel0),    //     conduit_control.export
		.channel1      (channel1),    //                    .export
		.fifo_status   (fifo_status), //                    .export
		.fifo_reset    (fifo_reset),  //                    .export
		.reg_address   (3'b000),      //         (terminated)
		.reg_write     (1'b0),        //         (terminated)
		.reg_writedata (8'b00000000), //         (terminated)
		.reg_read      (1'b0),        //         (terminated)
		.reg_readdata  ()             //         (terminated)
	);

endmodule
